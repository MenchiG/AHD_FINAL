----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:00:27 10/17/2016 
-- Design Name: 
-- Module Name:    ROM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ROM is
    Port ( address_i : in  STD_LOGIC_VECTOR (31 downto 0);
           data_o : out  STD_LOGIC_VECTOR (31 downto 0));
end ROM;

architecture Behavioral of ROM is

Type InstrMemType is array(natural range<>) of std_logic_vector(7 downto 0);  

constant Instruction : InstrMemtype:= (	  
"00011100","00000001","00000000","01101000", --0 a
"00011100","00000010","00000000","01101100", --4 b
"00011100","00000101","00000000","00000000", --8 s[0]
"00011100","00000100","00000000","00000100", --12 s[1]  
"00000000","00100011","00001000","00010000", --16 a+s[0]
"00000000","00100100","00001000","00010000", --20 b+s[1]
"00011100","00000100","00000000","01110100", --24 i<12
"00011100","00000101","00000000","01110000", --28 i=1
"00000000","00000001","00110000","00010100", --32 !a
"00000000","00000010","00111000","00010100", --36 !b
"00000000","11000010","01000000","00010010", --40
"00000000","11100001","01001000","00010010", --44
"00000001","00001001","01010000","00010011", --48 a xor b
"00001100","01001100","00000000","00011111", --52 j=amount
"00101000","00001100","00000000","00001100", --56 j==0? 
"00010101","01001010","00000000","00000001", --60 <<1
"00001001","10001100","00000000","00000001", --64 j--
"00101101","10000000","11111111","11110100", --68 j==0?
"00010100","10101101","00000000","00000011", --72 i*2*4
"00011101","10101110","00000000","00000000", --76 s[i*2*4]
"00000001","01001110","00001000","00010000", --80 a1
"00000000","00000001","00110000","00010100", --84 !a
"00000000","00000010","00111000","00010100", --88 !b
"00000000","11000010","01000000","00010010", --92
"00000000","11100001","01001000","00010010", --96
"00000001","00001001","01010000","00010011", --100 b xor a
"00001100","00101100","00000000","00011111", --104 j=amount
"00101000","00001100","00000000","00001100", --108 j==0? 
"00010101","01001010","00000000","00000001", --112 <<1
"00001001","10001100","00000000","00000001", --116 j--
"00101100","00001100","11111111","11110100", --120 j==0?
"00011101","10101110","00000000","00000100", --124 s[i*2*4+4]
"00000001","01001110","00010000","00010000", --128 b1
"00000100","10100101","00000000","00000001", --132 i++
"00101100","10000101","11111111","10010100", --136
"11111111","11111111","11111111","11111111"
);
begin


	 data_o <= Instruction(conv_integer(address_i)) & Instruction(conv_integer(address_i) + 1) & Instruction(conv_integer(address_i) + 2) & Instruction(conv_integer(address_i) + 3);
	 
end Behavioral;

